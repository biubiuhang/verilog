/* 3-8译码器设计

   abc              out
   000           0000_0001
   001           0000_0010
   010           0000_0100
   011           0000_1000
   100           0001_0000   
   101           0010_0000
   110           0100_0000
   111           1000_0000

*/

module decoder38(
   input        wire             a,
   input        wire             b,
   input        wire             c,
   output       reg    [7:0]     out
);

// 以always块描述的信号赋值，被赋值对象必须定义为reg类型

always@(*)
   case({a,b,c})
      3'b000:out = 8'b0000_0001;
      3'b001:out = 8'b0000_0010;
      3'b010:out = 8'b0000_0100;
      3'b011:out = 8'b0000_1000;
      3'b100:out = 8'b0001_0000;
      3'b101:out = 8'b0010_0000;
      3'b110:out = 8'b0100_0000;
      3'b111:out = 8'b1000_0000;
   endcase

// （{a,b,c}）变成一个三位的信号，这种操作叫做位拼接







endmodule
