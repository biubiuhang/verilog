/*
    时序逻辑基本概念（相较于之前的三八译码器）
    计数器基本概念，基本的4为加法器结构图
    设计一个以1s频率闪烁的LED灯（亮灭500ms）
    计数值与计数时间的关系
*/
module conter(
    input   wire              clk,
    input   wire              d,
    



); 








endmoudule